magic
tech scmos
timestamp 1699289289
<< nwell >>
rect -4 -16 314 66
<< ntransistor >>
rect 45 -37 53 -31
rect 114 -36 134 -32
rect 174 -36 194 -32
rect 242 -36 262 -32
rect 114 -67 134 -63
rect 169 -67 199 -63
rect 242 -67 262 -63
<< ptransistor >>
rect 214 28 290 33
rect 8 -2 90 2
rect 100 -2 148 2
rect 164 -5 204 5
rect 228 -2 276 2
<< ndiffusion >>
rect 45 -31 53 -30
rect 114 -30 120 -26
rect 128 -30 134 -26
rect 114 -32 134 -30
rect 174 -30 180 -26
rect 188 -30 194 -26
rect 174 -32 194 -30
rect 242 -30 248 -26
rect 256 -30 262 -26
rect 242 -32 262 -30
rect 45 -38 53 -37
rect 114 -38 134 -36
rect 114 -42 120 -38
rect 128 -42 134 -38
rect 174 -38 194 -36
rect 174 -42 180 -38
rect 188 -42 194 -38
rect 242 -38 262 -36
rect 242 -42 248 -38
rect 256 -42 262 -38
rect 114 -62 120 -58
rect 128 -62 134 -58
rect 114 -63 134 -62
rect 169 -62 180 -58
rect 188 -62 199 -58
rect 169 -63 199 -62
rect 242 -62 248 -58
rect 256 -62 262 -58
rect 242 -63 262 -62
rect 114 -68 134 -67
rect 114 -72 120 -68
rect 128 -72 134 -68
rect 169 -68 199 -67
rect 169 -72 180 -68
rect 188 -72 199 -68
rect 242 -68 262 -67
rect 242 -72 248 -68
rect 256 -72 262 -68
<< pdiffusion >>
rect 214 34 248 38
rect 256 34 290 38
rect 214 33 290 34
rect 214 27 290 28
rect 214 23 248 27
rect 256 23 290 27
rect 8 6 45 10
rect 53 6 90 10
rect 8 2 90 6
rect 100 6 120 10
rect 128 6 148 10
rect 100 2 148 6
rect 164 6 180 10
rect 188 6 204 10
rect 164 5 204 6
rect 228 6 248 10
rect 256 6 276 10
rect 8 -6 90 -2
rect 8 -10 45 -6
rect 53 -10 90 -6
rect 100 -6 148 -2
rect 228 2 276 6
rect 100 -10 120 -6
rect 128 -10 148 -6
rect 164 -6 204 -5
rect 164 -10 180 -6
rect 188 -10 204 -6
rect 228 -6 276 -2
rect 228 -10 248 -6
rect 256 -10 276 -6
<< ndcontact >>
rect 45 -30 53 -26
rect 120 -30 128 -26
rect 180 -30 188 -26
rect 248 -30 256 -26
rect 45 -42 53 -38
rect 120 -42 128 -38
rect 180 -42 188 -38
rect 248 -42 256 -38
rect 120 -62 128 -58
rect 180 -62 188 -58
rect 248 -62 256 -58
rect 120 -72 128 -68
rect 180 -72 188 -68
rect 248 -72 256 -68
<< pdcontact >>
rect 248 34 256 38
rect 248 23 256 27
rect 45 6 53 10
rect 120 6 128 10
rect 180 6 188 10
rect 248 6 256 10
rect 45 -10 53 -6
rect 120 -10 128 -6
rect 180 -10 188 -6
rect 248 -10 256 -6
<< psubstratepcontact >>
rect 0 -96 8 -88
rect 22 -96 30 -88
rect 45 -96 53 -88
rect 79 -96 95 -88
rect 120 -96 128 -88
rect 146 -96 162 -88
rect 180 -96 188 -88
rect 210 -96 226 -88
rect 248 -96 256 -88
rect 270 -96 278 -88
rect 290 -96 298 -88
<< nsubstratencontact >>
rect 0 54 8 62
rect 22 54 30 62
rect 45 54 53 62
rect 81 54 97 62
rect 120 54 128 62
rect 146 54 162 62
rect 180 54 188 62
rect 211 54 227 62
rect 248 54 256 62
rect 270 54 278 62
rect 290 54 298 62
<< polysilicon >>
rect 210 28 214 33
rect 290 28 294 33
rect 298 28 310 33
rect 0 -2 8 2
rect 148 -2 152 2
rect 160 -5 164 5
rect 204 -5 208 5
rect 212 -2 228 2
rect 276 -2 310 2
rect 41 -37 45 -31
rect 53 -32 57 -31
rect 53 -36 70 -32
rect 74 -36 114 -32
rect 134 -36 174 -32
rect 194 -36 242 -32
rect 262 -36 310 -32
rect 53 -37 57 -36
rect 110 -67 114 -63
rect 134 -67 144 -63
rect 148 -67 169 -63
rect 199 -67 242 -63
rect 262 -67 266 -63
<< polycontact >>
rect 294 28 298 33
rect 208 -5 212 5
rect 70 -36 74 -32
rect 144 -67 148 -63
<< polypplus >>
rect 90 -2 100 2
<< metal1 >>
rect 8 54 22 62
rect 30 54 45 62
rect 53 54 81 62
rect 97 54 120 62
rect 128 54 146 62
rect 162 54 180 62
rect 188 54 211 62
rect 227 54 248 62
rect 256 54 270 62
rect 278 54 290 62
rect 45 10 53 54
rect 120 10 128 54
rect 180 10 188 54
rect 248 38 256 54
rect 248 10 256 23
rect 45 -18 53 -10
rect 120 -18 128 -10
rect 180 -18 188 -10
rect 208 -18 212 -5
rect 45 -22 74 -18
rect 45 -26 53 -22
rect 70 -32 74 -22
rect 120 -22 148 -18
rect 120 -26 128 -22
rect 45 -88 53 -42
rect 120 -58 128 -42
rect 144 -63 148 -22
rect 180 -22 212 -18
rect 248 -18 256 -10
rect 294 -18 298 28
rect 248 -22 298 -18
rect 180 -26 188 -22
rect 248 -26 256 -22
rect 180 -58 188 -42
rect 248 -58 256 -42
rect 120 -88 128 -72
rect 180 -88 188 -72
rect 248 -88 256 -72
rect 8 -96 22 -88
rect 30 -96 45 -88
rect 53 -96 79 -88
rect 95 -96 120 -88
rect 128 -96 146 -88
rect 162 -96 180 -88
rect 188 -96 210 -88
rect 226 -96 248 -88
rect 256 -96 270 -88
rect 278 -96 290 -88
<< labels >>
rlabel polysilicon 0 -2 0 2 3 Vbias
rlabel polysilicon 310 28 310 33 7 Vbias4
rlabel polysilicon 310 -2 310 2 7 Vbias3
rlabel polysilicon 310 -36 310 -32 7 Vbias2
rlabel metal1 66 -92 66 -92 1 gnd!
rlabel metal1 66 58 66 58 1 Vdd!
<< end >>
